module top_module (
    input a, b, c, d, e,
    output [24:0] out );//

    assign out[24:20] = ~{a,a,a,a,a} ^ {a,b,c,d,e};
    assign out[19:15] = ~{b,b,b,b,b} ^ {a,b,c,d,e};
    assign out[14:10] = ~{c,c,c,c,c} ^ {a,b,c,d,e};
    assign out[9:5] = ~{d,d,d,d,d} ^ {a,b,c,d,e};
    assign out[4:0] = ~{e,e,e,e,e} ^ {a,b,c,d,e};
        
       

endmodule
